module trabalho3(
	input k = 1,
   input l = 0,
	input CLOCK_50;
	output reset = 0,
	output s = x;
);
	always @ (poseger CLOCK_50);
	 if (reset);
		
	
	for x (k, l + 20);
		
		if () begin;
			k = k + 1
		end	
			
		else begin;

		end


			for n ;
			
				if() begin;
					l = l + 1
					
				end
				
				else begin;
				
				end
end
endmodule
